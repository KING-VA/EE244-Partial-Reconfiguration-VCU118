`ifndef GARNET_CONFIG_SVH
`define GARNET_CONFIG_SVH

`define PARTITION_MODULE example
// `undef DISABLE_DDRA
// `undef DISABLE_DDRB
// `undef DISABLE_DEBUG_BRIDGE

`endif
